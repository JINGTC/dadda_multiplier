module dadda_24_tb();
       reg [23:0] A;
		 reg [23:0] B;
		 wire [46:0]mul_result;
		 
		 dadda_24 U1(
		 .B(B),
		 .A(A),
		 .mul_result(mul_result)
		 );
		 
		 initial
		 begin
		 #0 
		 A=24'b000011101001010100000000;
		 B=24'b000001001101001000000000;
		 #10
		 A=24'b000000111110100000000000;
		 B=24'b000000111110100100000000;
		 #10
		 A=24'b000001111101000000000000;
		 B=24'b000001111101000100000000;
		 #10
		 A=24'b000010111011100000000000;
		 B=24'b000010111011100100000000;
		 #10 $finish;
		 end
		 
		 endmodule
		 